module minimized_module (
    input x0,
    output reg f
);

    always @(*) begin
        f = 1'b1;
    end

endmodule
